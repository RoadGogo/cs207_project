module key_filter_module(
	clk,              // ������������ʱ��: 50Mhz
	rst_n,            // �����������븴λ����
	key_in,           // ���밴���ź�
	flag_key           // ���һ��ʱ�ӵĸߵ�ƽ
);

localparam n = 5;//�����ĸ���

//===========================================================================
// PORT declarations
//===========================================================================						
input        clk; 
input        rst_n;
input  [n-1:0] key_in;
output [n-1:0] flag_key;

//�Ĵ�������
reg [21:0] count;
reg [n-1:0] key_scan; //����ɨ��ֵKEY

//===========================================================================
// ��������ֵ��20msɨ��һ��,����Ƶ��С�ڰ���ë��Ƶ�ʣ��൱���˳����˸�Ƶë���źš�
//===========================================================================
always @(posedge clk or negedge rst_n)     //���ʱ�ӵ������غ͸�λ���½���
begin
   if(!rst_n)                //��λ�źŵ���Ч
	begin
      count <= 22'd0;        //��������0
		key_scan <= 0;
	end
   else
      begin
         if(count ==22'd1999_999)   //20msɨ��һ�ΰ���,20ms����(100M/50-1=1999_999)
         //if(count ==22'd2)//�����ڷ�����
            begin
               count <= 22'd0;     //�������Ƶ�20ms������������
               key_scan <= key_in; //�������������ƽ
            end
         else
            count <= count + 22'd1; //��������1
     end
end
//===========================================================================
// �����ź�����һ��ʱ�ӽ���
//===========================================================================
reg [n-1:0] key_scan_r = 0;
always @(posedge clk)
    key_scan_r <= key_scan;       
    
assign flag_key = key_scan_r[n-1:0] & (~key_scan[n-1:0]);  //����⵽�������Ͻ��ر仯ʱ������ð��������£�������Ч 

endmodule
